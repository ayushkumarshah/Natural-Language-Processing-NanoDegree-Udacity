BZh91AY&SY�`N _�Py���߰?���`��@��PJ�J$sFLL LFi�#ɀFѓ �`A��2`�4d���`F�b0L�a�101��&"�	��y�D	��F�4CF�=@�A4SBS�M�S�f�j��C�~�G���Q@{j,��8�R�J�	�x��K#��L�Q��g�c���EG�(\`��9@}��]М�[�#ƖA��M�% ��FQ|����@4�Z�:'��z$��			}5�L�1u�&���A(�$�ԧJ��fT�*x�t�c:F4�C�:�D�X� �5��v�Cg ,'$�����;�7֝�5��4�'�,�Jw�JY)��n��f�꣼��"%��ZE��<�.f�g���X�P�E�aX�$JN�>��F�5���H�5��p��g7Yn�f�I$�I��,E��:�8��8�C8�2�f	��zҫ�a4.P{�(���i�:
���F��82%l���� �~�OА��FH2I$�Jy'�|@�F#͉#�{@�ep,��Y=���%��L�g�B(���V�R%i��MhHHZ�P� 5���&͆�8	�tBA3����8}ծ/�1��>�g�:�<������u!3��u=�pJ)��3��|S�߀f�Ė����IPd�:�3B�Pzx�cw�����螴����Iަ;�P�'0��`i���j�q%Ɂ(~�*T���@�@�^@C}3��M�7�)�żHh� �`2��GJ�
�%�P���DB�n?�{'؝��h�^����1�8�6	�iJ��55�Z=olV���q5�� %�;%���*��	D�bPj��҂\��A��O�j@��t�~���B'�5P�D�\��H�8Z����T�Or���y�؇�@����DrD��it��⥉vdҍ���(���R�	��o��&5ʎ��m\jbxs�e���= ��8*�I�>�4�L`5�ɻ
'*t"@��p��M��
����- �2A��)�O��ĳB��D��pu�T���*#`"f��0�`�-�n�ː��NH�+U">�Z�m-ZlJ�c{ 0h�����ԚƆ�}#�p��	��'K�x@t�ArPe��ʗ7��� zUM��L�鼑��'4�(��C���'�ڝj��|��<�S��!��㰁��"H�%+P��qf ��i,&��R�����t��.�n��[�]2J��m=�u)�J%A�f�'SB��p��B�OY�Xz��P�ܛ n=��"��%C�<� ?I̛�b3���p9oC �c\*:������%�0�U�j�M�3�.�p�!����